`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Jafet Andr�s Chaves Barrantes
// 
// Create Date:    15:16:17 02/21/2016 
// Design Name: 
// Module Name:    Frecuency_Divider 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Frecuency_Divider(
    );


endmodule
